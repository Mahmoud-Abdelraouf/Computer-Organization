library verilog;
use verilog.vl_types.all;
entity PriorityResolver_tbFixedPriorities is
end PriorityResolver_tbFixedPriorities;
