library verilog;
use verilog.vl_types.all;
entity PriorityResolver_tbAutoRotation is
end PriorityResolver_tbAutoRotation;
