
module PriorityResolver_tb();
  
  
  
  
endmodule