library verilog;
use verilog.vl_types.all;
entity PriorityResolver_tb is
end PriorityResolver_tb;
