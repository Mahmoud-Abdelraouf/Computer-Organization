module RegisterFile (
    ports
);
    
endmodule