library verilog;
use verilog.vl_types.all;
entity InterruptMaskRegister_tb is
end InterruptMaskRegister_tb;
